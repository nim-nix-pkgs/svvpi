// Time-stamp: <2021-05-13 21:01:49 kmodi>

program top;

  initial begin
    $hello;
    $bye;
    void'($do_nothing);
    $finish;
  end

endprogram : top
